/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

module table_lookup (clk, state, p0, p1, p2, p3);
    input clk;
    input [31:0] state;
    output [31:0] p0, p1, p2, p3;
    wire [7:0] b0, b1, b2, b3;
    
    assign {b0, b1, b2, b3} = state;
    T
        t0 (clk, b0, {p0[23:0], p0[31:24]}),
        t1 (clk, b1, {p1[15:0], p1[31:16]}),
        t2 (clk, b2, {p2[7:0],  p2[31:8]} ),
        t3 (clk, b3, p3);
endmodule

/* substitue four bytes in a word */
module S4 (clk, in, out);
    input clk;
    input [31:0] in;
    output [31:0] out;
    
    S
        S_0 (clk, in[31:24], out[31:24]),
        S_1 (clk, in[23:16], out[23:16]),
        S_2 (clk, in[15:8],  out[15:8] ),
        S_3 (clk, in[7:0],   out[7:0]  );
endmodule

/* S_box, S_box, S_box*(x+1), S_box*x */
module T (clk, in, out);
    input clk;
    input [7:0] in;
    output reg [31:0] out;
    
    always @ (posedge clk)
    case (in)
    8'h00: out <= 32'h6363a5c6;
    8'h01: out <= 32'h7c7c84f8;
    8'h02: out <= 32'h777799ee;
    8'h03: out <= 32'h7b7b8df6;
    8'h04: out <= 32'hf2f20dff;
    8'h05: out <= 32'h6b6bbdd6;
    8'h06: out <= 32'h6f6fb1de;
    8'h07: out <= 32'hc5c55491;
    8'h08: out <= 32'h30305060;
    8'h09: out <= 32'h01010302;
    8'h0a: out <= 32'h6767a9ce;
    8'h0b: out <= 32'h2b2b7d56;
    8'h0c: out <= 32'hfefe19e7;
    8'h0d: out <= 32'hd7d762b5;
    8'h0e: out <= 32'hababe64d;
    8'h0f: out <= 32'h76769aec;
    8'h10: out <= 32'hcaca458f;
    8'h11: out <= 32'h82829d1f;
    8'h12: out <= 32'hc9c94089;
    8'h13: out <= 32'h7d7d87fa;
    8'h14: out <= 32'hfafa15ef;
    8'h15: out <= 32'h5959ebb2;
    8'h16: out <= 32'h4747c98e;
    8'h17: out <= 32'hf0f00bfb;
    8'h18: out <= 32'hadadec41;
    8'h19: out <= 32'hd4d467b3;
    8'h1a: out <= 32'ha2a2fd5f;
    8'h1b: out <= 32'hafafea45;
    8'h1c: out <= 32'h9c9cbf23;
    8'h1d: out <= 32'ha4a4f753;
    8'h1e: out <= 32'h727296e4;
    8'h1f: out <= 32'hc0c05b9b;
    8'h20: out <= 32'hb7b7c275;
    8'h21: out <= 32'hfdfd1ce1;
    8'h22: out <= 32'h9393ae3d;
    8'h23: out <= 32'h26266a4c;
    8'h24: out <= 32'h36365a6c;
    8'h25: out <= 32'h3f3f417e;
    8'h26: out <= 32'hf7f702f5;
    8'h27: out <= 32'hcccc4f83;
    8'h28: out <= 32'h34345c68;
    8'h29: out <= 32'ha5a5f451;
    8'h2a: out <= 32'he5e534d1;
    8'h2b: out <= 32'hf1f108f9;
    8'h2c: out <= 32'h717193e2;
    8'h2d: out <= 32'hd8d873ab;
    8'h2e: out <= 32'h31315362;
    8'h2f: out <= 32'h15153f2a;
    8'h30: out <= 32'h04040c08;
    8'h31: out <= 32'hc7c75295;
    8'h32: out <= 32'h23236546;
    8'h33: out <= 32'hc3c35e9d;
    8'h34: out <= 32'h18182830;
    8'h35: out <= 32'h9696a137;
    8'h36: out <= 32'h05050f0a;
    8'h37: out <= 32'h9a9ab52f;
    8'h38: out <= 32'h0707090e;
    8'h39: out <= 32'h12123624;
    8'h3a: out <= 32'h80809b1b;
    8'h3b: out <= 32'he2e23ddf;
    8'h3c: out <= 32'hebeb26cd;
    8'h3d: out <= 32'h2727694e;
    8'h3e: out <= 32'hb2b2cd7f;
    8'h3f: out <= 32'h75759fea;
    8'h40: out <= 32'h09091b12;
    8'h41: out <= 32'h83839e1d;
    8'h42: out <= 32'h2c2c7458;
    8'h43: out <= 32'h1a1a2e34;
    8'h44: out <= 32'h1b1b2d36;
    8'h45: out <= 32'h6e6eb2dc;
    8'h46: out <= 32'h5a5aeeb4;
    8'h47: out <= 32'ha0a0fb5b;
    8'h48: out <= 32'h5252f6a4;
    8'h49: out <= 32'h3b3b4d76;
    8'h4a: out <= 32'hd6d661b7;
    8'h4b: out <= 32'hb3b3ce7d;
    8'h4c: out <= 32'h29297b52;
    8'h4d: out <= 32'he3e33edd;
    8'h4e: out <= 32'h2f2f715e;
    8'h4f: out <= 32'h84849713;
    8'h50: out <= 32'h5353f5a6;
    8'h51: out <= 32'hd1d168b9;
    8'h52: out <= 32'h00000000;
    8'h53: out <= 32'heded2cc1;
    8'h54: out <= 32'h20206040;
    8'h55: out <= 32'hfcfc1fe3;
    8'h56: out <= 32'hb1b1c879;
    8'h57: out <= 32'h5b5bedb6;
    8'h58: out <= 32'h6a6abed4;
    8'h59: out <= 32'hcbcb468d;
    8'h5a: out <= 32'hbebed967;
    8'h5b: out <= 32'h39394b72;
    8'h5c: out <= 32'h4a4ade94;
    8'h5d: out <= 32'h4c4cd498;
    8'h5e: out <= 32'h5858e8b0;
    8'h5f: out <= 32'hcfcf4a85;
    8'h60: out <= 32'hd0d06bbb;
    8'h61: out <= 32'hefef2ac5;
    8'h62: out <= 32'haaaae54f;
    8'h63: out <= 32'hfbfb16ed;
    8'h64: out <= 32'h4343c586;
    8'h65: out <= 32'h4d4dd79a;
    8'h66: out <= 32'h33335566;
    8'h67: out <= 32'h85859411;
    8'h68: out <= 32'h4545cf8a;
    8'h69: out <= 32'hf9f910e9;
    8'h6a: out <= 32'h02020604;
    8'h6b: out <= 32'h7f7f81fe;
    8'h6c: out <= 32'h5050f0a0;
    8'h6d: out <= 32'h3c3c4478;
    8'h6e: out <= 32'h9f9fba25;
    8'h6f: out <= 32'ha8a8e34b;
    8'h70: out <= 32'h5151f3a2;
    8'h71: out <= 32'ha3a3fe5d;
    8'h72: out <= 32'h4040c080;
    8'h73: out <= 32'h8f8f8a05;
    8'h74: out <= 32'h9292ad3f;
    8'h75: out <= 32'h9d9dbc21;
    8'h76: out <= 32'h38384870;
    8'h77: out <= 32'hf5f504f1;
    8'h78: out <= 32'hbcbcdf63;
    8'h79: out <= 32'hb6b6c177;
    8'h7a: out <= 32'hdada75af;
    8'h7b: out <= 32'h21216342;
    8'h7c: out <= 32'h10103020;
    8'h7d: out <= 32'hffff1ae5;
    8'h7e: out <= 32'hf3f30efd;
    8'h7f: out <= 32'hd2d26dbf;
    8'h80: out <= 32'hcdcd4c81;
    8'h81: out <= 32'h0c0c1418;
    8'h82: out <= 32'h13133526;
    8'h83: out <= 32'hecec2fc3;
    8'h84: out <= 32'h5f5fe1be;
    8'h85: out <= 32'h9797a235;
    8'h86: out <= 32'h4444cc88;
    8'h87: out <= 32'h1717392e;
    8'h88: out <= 32'hc4c45793;
    8'h89: out <= 32'ha7a7f255;
    8'h8a: out <= 32'h7e7e82fc;
    8'h8b: out <= 32'h3d3d477a;
    8'h8c: out <= 32'h6464acc8;
    8'h8d: out <= 32'h5d5de7ba;
    8'h8e: out <= 32'h19192b32;
    8'h8f: out <= 32'h737395e6;
    8'h90: out <= 32'h6060a0c0;
    8'h91: out <= 32'h81819819;
    8'h92: out <= 32'h4f4fd19e;
    8'h93: out <= 32'hdcdc7fa3;
    8'h94: out <= 32'h22226644;
    8'h95: out <= 32'h2a2a7e54;
    8'h96: out <= 32'h9090ab3b;
    8'h97: out <= 32'h8888830b;
    8'h98: out <= 32'h4646ca8c;
    8'h99: out <= 32'heeee29c7;
    8'h9a: out <= 32'hb8b8d36b;
    8'h9b: out <= 32'h14143c28;
    8'h9c: out <= 32'hdede79a7;
    8'h9d: out <= 32'h5e5ee2bc;
    8'h9e: out <= 32'h0b0b1d16;
    8'h9f: out <= 32'hdbdb76ad;
    8'ha0: out <= 32'he0e03bdb;
    8'ha1: out <= 32'h32325664;
    8'ha2: out <= 32'h3a3a4e74;
    8'ha3: out <= 32'h0a0a1e14;
    8'ha4: out <= 32'h4949db92;
    8'ha5: out <= 32'h06060a0c;
    8'ha6: out <= 32'h24246c48;
    8'ha7: out <= 32'h5c5ce4b8;
    8'ha8: out <= 32'hc2c25d9f;
    8'ha9: out <= 32'hd3d36ebd;
    8'haa: out <= 32'hacacef43;
    8'hab: out <= 32'h6262a6c4;
    8'hac: out <= 32'h9191a839;
    8'had: out <= 32'h9595a431;
    8'hae: out <= 32'he4e437d3;
    8'haf: out <= 32'h79798bf2;
    8'hb0: out <= 32'he7e732d5;
    8'hb1: out <= 32'hc8c8438b;
    8'hb2: out <= 32'h3737596e;
    8'hb3: out <= 32'h6d6db7da;
    8'hb4: out <= 32'h8d8d8c01;
    8'hb5: out <= 32'hd5d564b1;
    8'hb6: out <= 32'h4e4ed29c;
    8'hb7: out <= 32'ha9a9e049;
    8'hb8: out <= 32'h6c6cb4d8;
    8'hb9: out <= 32'h5656faac;
    8'hba: out <= 32'hf4f407f3;
    8'hbb: out <= 32'heaea25cf;
    8'hbc: out <= 32'h6565afca;
    8'hbd: out <= 32'h7a7a8ef4;
    8'hbe: out <= 32'haeaee947;
    8'hbf: out <= 32'h08081810;
    8'hc0: out <= 32'hbabad56f;
    8'hc1: out <= 32'h787888f0;
    8'hc2: out <= 32'h25256f4a;
    8'hc3: out <= 32'h2e2e725c;
    8'hc4: out <= 32'h1c1c2438;
    8'hc5: out <= 32'ha6a6f157;
    8'hc6: out <= 32'hb4b4c773;
    8'hc7: out <= 32'hc6c65197;
    8'hc8: out <= 32'he8e823cb;
    8'hc9: out <= 32'hdddd7ca1;
    8'hca: out <= 32'h74749ce8;
    8'hcb: out <= 32'h1f1f213e;
    8'hcc: out <= 32'h4b4bdd96;
    8'hcd: out <= 32'hbdbddc61;
    8'hce: out <= 32'h8b8b860d;
    8'hcf: out <= 32'h8a8a850f;
    8'hd0: out <= 32'h707090e0;
    8'hd1: out <= 32'h3e3e427c;
    8'hd2: out <= 32'hb5b5c471;
    8'hd3: out <= 32'h6666aacc;
    8'hd4: out <= 32'h4848d890;
    8'hd5: out <= 32'h03030506;
    8'hd6: out <= 32'hf6f601f7;
    8'hd7: out <= 32'h0e0e121c;
    8'hd8: out <= 32'h6161a3c2;
    8'hd9: out <= 32'h35355f6a;
    8'hda: out <= 32'h5757f9ae;
    8'hdb: out <= 32'hb9b9d069;
    8'hdc: out <= 32'h86869117;
    8'hdd: out <= 32'hc1c15899;
    8'hde: out <= 32'h1d1d273a;
    8'hdf: out <= 32'h9e9eb927;
    8'he0: out <= 32'he1e138d9;
    8'he1: out <= 32'hf8f813eb;
    8'he2: out <= 32'h9898b32b;
    8'he3: out <= 32'h11113322;
    8'he4: out <= 32'h6969bbd2;
    8'he5: out <= 32'hd9d970a9;
    8'he6: out <= 32'h8e8e8907;
    8'he7: out <= 32'h9494a733;
    8'he8: out <= 32'h9b9bb62d;
    8'he9: out <= 32'h1e1e223c;
    8'hea: out <= 32'h87879215;
    8'heb: out <= 32'he9e920c9;
    8'hec: out <= 32'hcece4987;
    8'hed: out <= 32'h5555ffaa;
    8'hee: out <= 32'h28287850;
    8'hef: out <= 32'hdfdf7aa5;
    8'hf0: out <= 32'h8c8c8f03;
    8'hf1: out <= 32'ha1a1f859;
    8'hf2: out <= 32'h89898009;
    8'hf3: out <= 32'h0d0d171a;
    8'hf4: out <= 32'hbfbfda65;
    8'hf5: out <= 32'he6e631d7;
    8'hf6: out <= 32'h4242c684;
    8'hf7: out <= 32'h6868b8d0;
    8'hf8: out <= 32'h4141c382;
    8'hf9: out <= 32'h9999b029;
    8'hfa: out <= 32'h2d2d775a;
    8'hfb: out <= 32'h0f0f111e;
    8'hfc: out <= 32'hb0b0cb7b;
    8'hfd: out <= 32'h5454fca8;
    8'hfe: out <= 32'hbbbbd66d;
    8'hff: out <= 32'h16163a2c;
    endcase
endmodule

/* S box */
module S (clk, in, out);
    input clk;
    input [7:0] in;
    output reg [7:0] out;

    always @ (posedge clk)
    case (in)
    8'h00: out <= 8'h63;
    8'h01: out <= 8'h7c;
    8'h02: out <= 8'h77;
    8'h03: out <= 8'h7b;
    8'h04: out <= 8'hf2;
    8'h05: out <= 8'h6b;
    8'h06: out <= 8'h6f;
    8'h07: out <= 8'hc5;
    8'h08: out <= 8'h30;
    8'h09: out <= 8'h01;
    8'h0a: out <= 8'h67;
    8'h0b: out <= 8'h2b;
    8'h0c: out <= 8'hfe;
    8'h0d: out <= 8'hd7;
    8'h0e: out <= 8'hab;
    8'h0f: out <= 8'h76;
    8'h10: out <= 8'hca;
    8'h11: out <= 8'h82;
    8'h12: out <= 8'hc9;
    8'h13: out <= 8'h7d;
    8'h14: out <= 8'hfa;
    8'h15: out <= 8'h59;
    8'h16: out <= 8'h47;
    8'h17: out <= 8'hf0;
    8'h18: out <= 8'had;
    8'h19: out <= 8'hd4;
    8'h1a: out <= 8'ha2;
    8'h1b: out <= 8'haf;
    8'h1c: out <= 8'h9c;
    8'h1d: out <= 8'ha4;
    8'h1e: out <= 8'h72;
    8'h1f: out <= 8'hc0;
    8'h20: out <= 8'hb7;
    8'h21: out <= 8'hfd;
    8'h22: out <= 8'h93;
    8'h23: out <= 8'h26;
    8'h24: out <= 8'h36;
    8'h25: out <= 8'h3f;
    8'h26: out <= 8'hf7;
    8'h27: out <= 8'hcc;
    8'h28: out <= 8'h34;
    8'h29: out <= 8'ha5;
    8'h2a: out <= 8'he5;
    8'h2b: out <= 8'hf1;
    8'h2c: out <= 8'h71;
    8'h2d: out <= 8'hd8;
    8'h2e: out <= 8'h31;
    8'h2f: out <= 8'h15;
    8'h30: out <= 8'h04;
    8'h31: out <= 8'hc7;
    8'h32: out <= 8'h23;
    8'h33: out <= 8'hc3;
    8'h34: out <= 8'h18;
    8'h35: out <= 8'h96;
    8'h36: out <= 8'h05;
    8'h37: out <= 8'h9a;
    8'h38: out <= 8'h07;
    8'h39: out <= 8'h12;
    8'h3a: out <= 8'h80;
    8'h3b: out <= 8'he2;
    8'h3c: out <= 8'heb;
    8'h3d: out <= 8'h27;
    8'h3e: out <= 8'hb2;
    8'h3f: out <= 8'h75;
    8'h40: out <= 8'h09;
    8'h41: out <= 8'h83;
    8'h42: out <= 8'h2c;
    8'h43: out <= 8'h1a;
    8'h44: out <= 8'h1b;
    8'h45: out <= 8'h6e;
    8'h46: out <= 8'h5a;
    8'h47: out <= 8'ha0;
    8'h48: out <= 8'h52;
    8'h49: out <= 8'h3b;
    8'h4a: out <= 8'hd6;
    8'h4b: out <= 8'hb3;
    8'h4c: out <= 8'h29;
    8'h4d: out <= 8'he3;
    8'h4e: out <= 8'h2f;
    8'h4f: out <= 8'h84;
    8'h50: out <= 8'h53;
    8'h51: out <= 8'hd1;
    8'h52: out <= 8'h00;
    8'h53: out <= 8'hed;
    8'h54: out <= 8'h20;
    8'h55: out <= 8'hfc;
    8'h56: out <= 8'hb1;
    8'h57: out <= 8'h5b;
    8'h58: out <= 8'h6a;
    8'h59: out <= 8'hcb;
    8'h5a: out <= 8'hbe;
    8'h5b: out <= 8'h39;
    8'h5c: out <= 8'h4a;
    8'h5d: out <= 8'h4c;
    8'h5e: out <= 8'h58;
    8'h5f: out <= 8'hcf;
    8'h60: out <= 8'hd0;
    8'h61: out <= 8'hef;
    8'h62: out <= 8'haa;
    8'h63: out <= 8'hfb;
    8'h64: out <= 8'h43;
    8'h65: out <= 8'h4d;
    8'h66: out <= 8'h33;
    8'h67: out <= 8'h85;
    8'h68: out <= 8'h45;
    8'h69: out <= 8'hf9;
    8'h6a: out <= 8'h02;
    8'h6b: out <= 8'h7f;
    8'h6c: out <= 8'h50;
    8'h6d: out <= 8'h3c;
    8'h6e: out <= 8'h9f;
    8'h6f: out <= 8'ha8;
    8'h70: out <= 8'h51;
    8'h71: out <= 8'ha3;
    8'h72: out <= 8'h40;
    8'h73: out <= 8'h8f;
    8'h74: out <= 8'h92;
    8'h75: out <= 8'h9d;
    8'h76: out <= 8'h38;
    8'h77: out <= 8'hf5;
    8'h78: out <= 8'hbc;
    8'h79: out <= 8'hb6;
    8'h7a: out <= 8'hda;
    8'h7b: out <= 8'h21;
    8'h7c: out <= 8'h10;
    8'h7d: out <= 8'hff;
    8'h7e: out <= 8'hf3;
    8'h7f: out <= 8'hd2;
    8'h80: out <= 8'hcd;
    8'h81: out <= 8'h0c;
    8'h82: out <= 8'h13;
    8'h83: out <= 8'hec;
    8'h84: out <= 8'h5f;
    8'h85: out <= 8'h97;
    8'h86: out <= 8'h44;
    8'h87: out <= 8'h17;
    8'h88: out <= 8'hc4;
    8'h89: out <= 8'ha7;
    8'h8a: out <= 8'h7e;
    8'h8b: out <= 8'h3d;
    8'h8c: out <= 8'h64;
    8'h8d: out <= 8'h5d;
    8'h8e: out <= 8'h19;
    8'h8f: out <= 8'h73;
    8'h90: out <= 8'h60;
    8'h91: out <= 8'h81;
    8'h92: out <= 8'h4f;
    8'h93: out <= 8'hdc;
    8'h94: out <= 8'h22;
    8'h95: out <= 8'h2a;
    8'h96: out <= 8'h90;
    8'h97: out <= 8'h88;
    8'h98: out <= 8'h46;
    8'h99: out <= 8'hee;
    8'h9a: out <= 8'hb8;
    8'h9b: out <= 8'h14;
    8'h9c: out <= 8'hde;
    8'h9d: out <= 8'h5e;
    8'h9e: out <= 8'h0b;
    8'h9f: out <= 8'hdb;
    8'ha0: out <= 8'he0;
    8'ha1: out <= 8'h32;
    8'ha2: out <= 8'h3a;
    8'ha3: out <= 8'h0a;
    8'ha4: out <= 8'h49;
    8'ha5: out <= 8'h06;
    8'ha6: out <= 8'h24;
    8'ha7: out <= 8'h5c;
    8'ha8: out <= 8'hc2;
    8'ha9: out <= 8'hd3;
    8'haa: out <= 8'hac;
    8'hab: out <= 8'h62;
    8'hac: out <= 8'h91;
    8'had: out <= 8'h95;
    8'hae: out <= 8'he4;
    8'haf: out <= 8'h79;
    8'hb0: out <= 8'he7;
    8'hb1: out <= 8'hc8;
    8'hb2: out <= 8'h37;
    8'hb3: out <= 8'h6d;
    8'hb4: out <= 8'h8d;
    8'hb5: out <= 8'hd5;
    8'hb6: out <= 8'h4e;
    8'hb7: out <= 8'ha9;
    8'hb8: out <= 8'h6c;
    8'hb9: out <= 8'h56;
    8'hba: out <= 8'hf4;
    8'hbb: out <= 8'hea;
    8'hbc: out <= 8'h65;
    8'hbd: out <= 8'h7a;
    8'hbe: out <= 8'hae;
    8'hbf: out <= 8'h08;
    8'hc0: out <= 8'hba;
    8'hc1: out <= 8'h78;
    8'hc2: out <= 8'h25;
    8'hc3: out <= 8'h2e;
    8'hc4: out <= 8'h1c;
    8'hc5: out <= 8'ha6;
    8'hc6: out <= 8'hb4;
    8'hc7: out <= 8'hc6;
    8'hc8: out <= 8'he8;
    8'hc9: out <= 8'hdd;
    8'hca: out <= 8'h74;
    8'hcb: out <= 8'h1f;
    8'hcc: out <= 8'h4b;
    8'hcd: out <= 8'hbd;
    8'hce: out <= 8'h8b;
    8'hcf: out <= 8'h8a;
    8'hd0: out <= 8'h70;
    8'hd1: out <= 8'h3e;
    8'hd2: out <= 8'hb5;
    8'hd3: out <= 8'h66;
    8'hd4: out <= 8'h48;
    8'hd5: out <= 8'h03;
    8'hd6: out <= 8'hf6;
    8'hd7: out <= 8'h0e;
    8'hd8: out <= 8'h61;
    8'hd9: out <= 8'h35;
    8'hda: out <= 8'h57;
    8'hdb: out <= 8'hb9;
    8'hdc: out <= 8'h86;
    8'hdd: out <= 8'hc1;
    8'hde: out <= 8'h1d;
    8'hdf: out <= 8'h9e;
    8'he0: out <= 8'he1;
    8'he1: out <= 8'hf8;
    8'he2: out <= 8'h98;
    8'he3: out <= 8'h11;
    8'he4: out <= 8'h69;
    8'he5: out <= 8'hd9;
    8'he6: out <= 8'h8e;
    8'he7: out <= 8'h94;
    8'he8: out <= 8'h9b;
    8'he9: out <= 8'h1e;
    8'hea: out <= 8'h87;
    8'heb: out <= 8'he9;
    8'hec: out <= 8'hce;
    8'hed: out <= 8'h55;
    8'hee: out <= 8'h28;
    8'hef: out <= 8'hdf;
    8'hf0: out <= 8'h8c;
    8'hf1: out <= 8'ha1;
    8'hf2: out <= 8'h89;
    8'hf3: out <= 8'h0d;
    8'hf4: out <= 8'hbf;
    8'hf5: out <= 8'he6;
    8'hf6: out <= 8'h42;
    8'hf7: out <= 8'h68;
    8'hf8: out <= 8'h41;
    8'hf9: out <= 8'h99;
    8'hfa: out <= 8'h2d;
    8'hfb: out <= 8'h0f;
    8'hfc: out <= 8'hb0;
    8'hfd: out <= 8'h54;
    8'hfe: out <= 8'hbb;
    8'hff: out <= 8'h16;
    endcase
endmodule
